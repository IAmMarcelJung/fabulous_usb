`ifndef MACROS_VH
`define MACROS_VH

`define MAX(a,b) ((a) > (b) ? (a) : (b))
`define MIN(a,b) ((a) < (b) ? (a) : (b))

`endif
